`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Create Date: 01/26/2025 11:53:46 PM
// Design Name: UARTLedSystem
// Module Name: UARTLedSystem
// Project Name: UARTLedSystem
// Target Devices: Basys3
// Tool Versions: 2023.2
// Description: The top level module for the UARTLedSystem project.
//////////////////////////////////////////////////////////////////////////////////


module UARTLedSystem (
    input  wire        Clk,
    input  wire        Reset,
    input  wire        SentUartData,
    input  wire [ 7:0] Sw,
    output wire        UARTTx,
    input  wire        UARTRx,
    output wire [15:0] Led
);
  // Add your code here

  // End or your code
endmodule
